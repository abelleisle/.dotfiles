Vim�UnDo� Xj���96��fo�eh��\ �\����ϕ�Y㳀   m                                   Z�`@    _�                      E        ����                                                                                                                                                                                                                                                                                                                            E           �           V        Z�`@     �   F   G   m   &     -- stimulus CLK   $  CLK <= not CLK after clk_period/2;         -- stimulus RST     stimulusRST: process     begin   (      RST <= '1';            -- at  0 ns         wait for clk_period/4;     (      RST <= '0';            -- at 25 ns         wait for clk_period/2;     D      RST <= ____;           -- at 75 ns, fill in the new RST value          wait;     end process;   	       -- stimulus SL     stimulusSL: process     begin   (      SL <= '1';             -- at  0 ns         wait for 125 ns;          E      SL <= ____;            -- at 125 ns, fill in the new SL value           wait;     end process;       -- stimulus SIN     stimulusSIN: process     begin   (      SIN <= '0';            -- at  0 ns         wait for 325 ns;          F      SIN <= ____;           -- at 325 ns, fill in the new SIN value           wait;     end process;       -- stimulus A, B, C, D        4  A <= ____;                 -- fill in A value        0  B <= ____;                 -- fill in B value    /  C <= ____;                 -- fill in C value   2  D <= ____;                 -- fill in D value   5��